`include "ALU_iface.sv"
`include "environment.sv"

module test (ALU_iface ifc);

  environment env = new(ifc);

  initial
  begin
    $timeformat(-9,0," ns" , 10);
    env.run();
  end

endmodule : test
